library ieee;
  use ieee.std_logic_1164.all;

package foo is

  type t_my is record
    a : std_logic;
    b : std_logic;
  end record t_my;

end package foo;
