library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

package pkg is

  subtype foo is std_logic_vector(3 downto 0);

end package pkg;
